`ifdef USE_MODULE_CLKDIV

module Gowin_CLKDIV (clkout, hclkin, resetn);

    output clkout;
    input hclkin;
    input resetn;

    wire gw_gnd;

    assign gw_gnd = 1'b0;

    CLKDIV clkdiv_inst (
               .CLKOUT(clkout),
               .HCLKIN(hclkin),
               .RESETN(resetn),
               .CALIB(gw_gnd)
           );

    defparam clkdiv_inst.DIV_MODE = "2";
    defparam clkdiv_inst.GSREN = "false";

endmodule

`endif
