//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.09 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Tue Feb 28 21:26:49 2023

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din);

    output [7:0] dout;
    input clk;
    input oce;
    input ce;
    input reset;
    input wre;
    input [10:0] ad;
    input [7:0] din;

    wire [23:0] sp_inst_0_dout_w;
    wire gw_gnd;

    assign gw_gnd = 1'b0;

    SP sp_inst_0 (
           .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
           .CLK(clk),
           .OCE(oce),
           .CE(ce),
           .RESET(reset),
           .WRE(wre),
           .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
           .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
           .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
       );

    defparam sp_inst_0.READ_MODE = 1'b0;
    defparam sp_inst_0.WRITE_MODE = 2'b00;
    defparam sp_inst_0.BIT_WIDTH = 8;
    defparam sp_inst_0.BLK_SEL = 3'b000;
    defparam sp_inst_0.RESET_MODE = "SYNC";

    defparam sp_inst_0.INIT_RAM_00 = 256'hFEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210; // 256-bit: 64 hex (2 hex -> 1 byte)


endmodule //Gowin_SP
